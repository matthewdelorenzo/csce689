
    always @(posedge clk) begin
        q <= d;
    end

endmodule
