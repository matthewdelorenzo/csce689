//Please finish designing the 64 bit multiplier module (multiplier_64) below.
//There are two 64 bit inputs (A and B) and a 128 bit output (product).
//The module should utilize the inputs (A and B) to determine the output product correctly in its implementation.
module multiplier_64(output [127:0] product, input [63:0] A, B);
	
	wire [63:0] pp0, pp1, pp2, pp3, pp4, pp5, pp6, pp7, pp8, pp9, pp10, pp11, pp12, pp13, pp14, pp15;
	wire [63:0] pp16, pp17, pp18, pp19, pp20, pp21, pp22, pp23, pp24, pp25, pp26, pp27, pp28, pp29, pp30, pp31;
	wire [63:0] pp32, pp33, pp34, pp35, pp36, pp37, pp38, pp39, pp40, pp41, pp42, pp43, pp44, pp45, pp46, pp47;
	wire [63:0] pp48, pp49, pp50, pp51, pp52, pp53, pp54, pp55, pp56, pp57, pp58, pp59, pp60, pp61, pp62, pp63;
	wire [127:0] product1;
	wire [127:0] product2;
	wire [127:0] product3;
	wire [127:0] product4;
	wire [127:0] product5;
	wire [127:0] product6;
	wire [127:0] product7;
	wire [127:0] product8;
	wire [127:0] product9;
	wire [127:0] product10;
	wire [127:0] product11;
	wire [127:0] product12;
	wire [127:0] product13;
	wire [127:0] product14;
	wire [127:0] product15;
	wire [127:0] product16;
	wire [127:0] product17;
	wire [127:0] product18;
	wire [127:0] product19;
	wire [127:0] product20;
	wire [127:0] product21;
	wire [127:0] product22;
	wire [127:0] product23;
	wire [127:0] product24;
	wire [127:0] product25;
	wire [127:0] product26;
	wire [127:0] product27;
	wire [127:0] product28;
	wire [127:0] product29;
	wire [127:0] product30;
	wire [127:0] product31;
	wire [127:0] product32;
	wire [127:0] product33;
	wire [127:0] product34;
	wire [127:0] product35;
	wire [127:0] product36;
	wire [127:0] product37;
	wire [127:0] product38;
	wire [127:0] product39;
	wire [127:0] product40;
	wire [127:0] product41;
	wire [127:0] product42;
	wire [127:0] product43;
	wire [127:0] product44;
	wire [127:0] product45;
	wire [127:0] product46;
	wire [127:0] product47;
	wire [127:0] product48;
	wire [127:0] product49;
	wire [127:0] product50;
	wire [127:0] product51;
	wire [127:0] product52;
	wire [127:0] product53;
	wire [127:0] product54;
	wire [127:0] product55;
	wire [127:0] product56;
	wire [127:0] product57;
	wire [127:0] product58;
	wire [127:0] product59;
	wire [127:0] product60;
	wire [127:0] product61;
	wire [127:0] product62;
	wire [127:0] product63;
	wire [127:0] product64;
	
	assign pp0 = A[0]? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
	assign pp1 = A[1]? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
	assign pp2 = A[2]? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
	assign pp3 = A[3]? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
	assign