// Build a 32-bit Galois LFSR with taps at bit positions 32, 22, 2, and 1.

// Hint: This is long enough that you'd want to use vectors, not 32 instantiations of DFFs.

module top_module(
    input clk,
    input reset,    // Active-high synchronous reset to 32'h1
    output [31:0] q
); 
    
    reg [31:0] q_next;
    
    always @(*) begin
        q_next = q[31]? {q[30:0], 1'b0} : q_next;
    end
    
    always @(posedge clk) begin
        if(reset)
            q <= 32'h1;
        else
            q <= q_next;
    end
    
endmodule