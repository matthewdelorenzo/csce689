//Please finish designing the 32 bit multiplier module (multiplier_32) below.
//There are two 32 bit inputs (A and B) and a 64 bit output (product).
//The module should utilize the inputs (A and B) to determine the output product correctly in its implementation.
module multiplier_32(output [63:0] product, input [31:0] A, B);
	assign pp0 = A[0]? B: 32'b00000000000000000000000000000000;
	assign pp1 = A[1]? B: 32'b00000000000000000000000000000000;
	assign pp2 = A[2]? B: 32'b00000000000000000000000000000000;
	assign pp3 = A[3]? B: 32'b00000000000000000000000000000000;
	assign pp4 = A[4]? B: 32'b00000000000000000000000000000000;
	assign pp5 = A[5]? B: 32'b00000000000000000000000000000000;
	assign pp6 = A[6]? B: 32'b00000000000000000000000000000000;
	assign pp7 = A[7]? B: 32'b00000000000000000000000000000000;
	assign pp8 = A[8]? B: 32'b00000000000000000000000000000000;
	assign pp9 = A[9]? B: 32'b00000000000000000000000000000000;
	assign pp10 = A[10]? B: 32'b00000000000000000000000000000000;
	assign pp11 = A[11]? B: 32'b00000000000000000000000000000000;
	assign pp12 = A[12]? B: 32'b00000000000000000000000000000000;
	assign pp13 = A[13]? B: 32'b00000000000000000000000000000000;
	assign pp14 = A[14]? B: 32'b00000000000000000000000000000000;
	assign pp15 = A[15]? B: 32'b00000000000000000000000000000000;
	assign pp16 = A[16]? B: 32'b00000000000000000000000000000000;
	assign pp17 = A[17]? B: 32'b00000000000000000000000000000000;
	assign pp18 = A[18]? B: 32'b00000000000000000000000000000000;
	assign pp19 = A[19]? B: 32'b00000000000000000000000000000000;
	assign pp20 = A[20]? B: 32'b00000000000000000000000000000000;
	assign pp21 = A[21]? B: 32'b00000000000000000000000000000000;
	assign pp22 = A[22]? B: 32'b00000000000000000000000000000000;
	assign pp23 = A[23]? B: 32'b00000000000000000000000000000000;
	assign pp24 = A[24]? B: 32'b00000000000000000000000000000000;
	assign pp25 = A[25]? B: 32'b00000000000000000000000000000000;
	assign pp26 = A[26]? B: 32'b00000000000000000000000000000000;
	assign pp27 = A[27]? B: 32'b00000000000000000000000000000000;
	assign pp28 = A[28]? B: 32'b00000000000000000000000000000000;
	assign pp29 = A[29]? B: 32'b00000000000000000000000000000000;
	assign pp30 = A[30]? B: 32'b00000000000000000000000000000000;
	assign pp31 = A[31]? B: 32'b00000000000000000000000000000000;
	assign product[0] = pp0[0];
	assign in1_1 = {pp0[1],pp0[0],pp0[0],pp0[0]};
	assign in1_2 = {pp1[0],pp1[0],pp1[0],pp1[0]};
	CLA4 CLA01(s1, c1, in1_1, in1_2);
	assign in2_1 = {pp2[1],pp2[0],pp2[0],pp2[0]};
	assign in2_2 = {pp3[0],pp3[0],pp3[0],pp3[0]};
	CLA4 CLA02(s2, c2, in2_1, in2_2);
	assign in3_1 = {s1[3],s1[2],s1[1],s1[0]};
	assign in3_2 = {s2[2],s2[1],s2[0],s2[3]};
	CLA4 CLA03(s3, c3, in3_1, in3_2);
	assign in4_1 = {pp4[1],pp4[0],pp4[0],pp4[0]};
	assign in4_2 = {pp5[0],pp5[0],pp5[0],pp5[0]};
	CLA4 CLA04(s4, c4, in4_1, in4_2);
	assign in5_1 = {s1[3],s1[2],s1[1],s1[0]