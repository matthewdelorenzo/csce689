// create one instance of module mod_a, then connect the module's three pins (in1, in2, and out) 
// to your top-level module's three ports (wires a, b, and out). 
//The module mod_a is provided for you — you must instantiate it.


//Hint: When connecting modules, only the ports on the module are important. 
// You do not need to know the code inside the module. 
// The code for module mod_a looks like this:

module top_module ( input a, input b, output out );
mod_a instance_name (
        .in1(a), 
        .in2(b), 
        .out(out)
    );
endmodule