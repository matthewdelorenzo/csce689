    
    assign {cout, sum} = a + b;

endmodule
