    mod_a instance1(.out(out), .in1(a), .in2(b));
endmodule
