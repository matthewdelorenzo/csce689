    
    assign out = (~b & c) | (a & c) | (a & ~c);

endmodule
