
    assign out = in[sel*4+3 -: 4]; // - and : should be put together
    
endmodule
