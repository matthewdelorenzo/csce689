//Please finish designing the 64 bit multiplier module (multiplier_64) below.
//There are two 64 bit inputs (A and B) and a 128 bit output (product).
//The module should utilize the inputs (A and B) to determine the output product correctly in its implementation.
module multiplier_64(output [127:0] product, input [63:0] A, B); 

//Please fill in the code for the multiplier_64 module.
//You may use the following variables in your code:
 //A, B, product
//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code:
 //adder_64

//You may use the following modules in your code: