    assign parity = ^ in[7:0];
endmodule
