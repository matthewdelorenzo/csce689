//Please finish designing the 16 bit multiplier module (multiplier_16) below.
//There are two 16 bit inputs (A and B) and a 32 bit output (product).
//The module should utilize the inputs (A and B) to determine the output product correctly in its implementation.
module top_module(output [31:0] product, input [15:0] A, B);

  assign product = A * B;
endmodule