//Please finish designing the 32 bit multiplier module (multiplier_32) below.
//There are two 32 bit inputs (A and B) and a 64 bit output (product).
//The module should utilize the inputs (A and B) to determine the output product correctly in its implementation.
module multiplier_32(output [63:0] product, input [31:0] A, B);

//Please finish implementing the 32 bit multiplier module (multiplier_32) below.
//There are two 32 bit inputs (A and B) and a 64 bit output (product).
//The module should utilize the inputs (A and B) to determine the output product correctly in its implementation.

//You may use any number of wires and logic gates to implement the multiplier.
//You may use the following 32 bit full adder module as a submodule in your implementation.
//The 32 bit full adder module is located in the following file:
//"C:\Users\johndoe\Desktop\School\ECE 341\Lab 2\full_adder_32.v"

//You may use the following 32 bit half adder module as a submodule in your implementation.
//The 32 bit half adder module is located in the following file:
//"C:\Users\johndoe\Desktop\School\ECE 341\Lab 2\half_adder_32.v"

//You may use the following 32 bit half adder module as a submodule in your implementation.
//The 32 bit half adder module is located in the following file:
//"C:\Users\johndoe\Desktop\School\ECE 341\Lab 2\half_adder_32.v"

//You may use the following 32 bit half adder module as a submodule in your implementation.
//The 32 bit half adder module is located in the following file:
//"C:\Users\johndoe\Desktop\School\ECE 341\Lab 2\half_adder_32.v"

//You may use the following 32 bit half adder module as a submodule in your implementation.
//The 32 bit half adder module is located in the following file:
//"C:\Users\johndoe\Desktop\School\ECE 341\Lab 2\half_adder_32.v"

//You may use the following 32 bit half adder module as a submodule in your implementation.
//The 32 bit half adder module is located in the following file:
//"C:\Users\johndoe\Desktop\School\ECE 341\Lab 2\half_adder_32.v"

//You may use the following 32 bit half adder module as a submodule in your implementation.
//The 32 bit half adder module is located in the following file:
//"C:\Users\johndoe\Desktop\School\ECE 341\Lab 2\half_adder_32.v"

//You may use the following 32 bit half adder module as a submodule in your implementation.
//The 32 bit half adder module is located in the following file:
//"C:\Users\johndoe\Desktop\School\ECE 341\Lab 2\half_adder_32.v"

//You may use the following 32 bit half adder module as a submodule in your implementation.
//The 32 bit half adder module is located in the following file:
//"C:\Users\johndoe\Desktop\School\ECE 341\Lab 2\half_adder_32.v"

//You may use the following 32 bit half adder module as a submodule in your implementation.
//The 32 bit half adder module is located in the following file:
//"C:\Users\johndoe\Desktop\School\ECE 341\Lab 2\half_adder_32.v"

//You may use the following 32 bit half adder module as a submodule in your implementation.
//The 32 bit half adder module is located in the following file:
//"C:\Users\johndoe\Desktop\School\ECE 341\Lab 2\half_adder_32.v"

//You may use the following 32 bit half adder module as a submodule in your implementation.
//The 32 bit half adder module is located in the following file:
//"C:\Users\johndoe\Desktop\School\ECE 341\Lab 2\half_adder_32.v"

//You may use the following 32 bit half adder module as a submodule in your implementation.
//The 32 bit half adder module is located in the following file:
//"C:\Users\johndoe\Desktop\School\ECE 341\Lab 2\half_adder_32.v"

//You may use the following 32 bit half adder module as a submodule in your implementation.
//The 32 bit half adder module is located in the following file:
//"C:\Users\johndoe\Desktop\School\ECE 341\Lab 2\half_adder_32.v"

//You may use the following 32 bit half adder module as a submodule in your implementation.
//The 32 bit half adder module is located in the following file:
//"C:\Users\johndoe\Desktop\School\ECE 341\Lab 2\half_adder_32.v"

//You may use the following 32 bit half adder module as a submodule in your implementation.
//The 32 bit half adder module is located in the following file:
//"C:\Users\johndoe\Desktop\School\ECE 341\Lab 2\half_adder_32.v"

//You may use the following 32 bit half adder module as a submodule in your implementation.
//The 32 bit half adder module is located in the following file:
//"C:\Users\johndoe\Desktop\School\ECE 341\Lab 2\half_adder_32.v"

//You may use the following 32 bit half adder module as a submodule in your implementation.
//The 32 bit half adder module is located in the following file:
//"C:\Users\johndoe\Desktop\School\ECE 341\Lab 2\half_adder_32.v"

//You may use the following 32 bit half adder module as a submodule in your implementation.
//The 32 bit half adder module is located in the following file:
//"C:\Users\johndoe\Desktop\School\ECE 341\Lab 2\half_adder_32.v"

//You may use the following 32 bit half adder module as a submodule in your implementation.
//The 32 bit half adder module is located in the following file:
//"C:\Users\johndoe\Desktop\School\ECE 341\Lab 2\half_adder_32.v"

//You may use the following 32 bit half adder module as a submodule in your implementation.
//The 32 bit half adder module is located in the following file:
//"C:\Users\johndoe\Desktop\School\ECE 341\Lab 2\half_adder_32.v"

//You may use the following 32 bit half adder module as a submodule in your implementation.
//The 32 bit half adder module is located in the following file:
//"C:\Users\johndoe\Desktop\School\ECE 341\Lab 2\half_adder_32.v"

//You may use the following 32 bit half adder module as a submodule in your implementation.
//The 32 bit half adder module is located in the following file:
//"C:\Users\johndoe\Desktop\School\ECE 341\Lab 2\half_adder_32.v"

//You may use the following 32 bit half adder module as a submodule in your implementation.
//The 32 bit half adder module is located in the following file:
//"C:\Users\johndoe\Desktop\School\ECE 341\Lab 2\half_adder_32.v"

//You may use the following 32 bit half adder module as a submodule in your implementation.
//The 32 bit half adder module is located in