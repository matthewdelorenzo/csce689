// You are provided with a BCD one-digit adder named bcd_fadd that adds 
// two BCD digits and carry-in, and produces a sum and carry-out.

module bcd_fadd (
    input [3:0] a,
    input [3:0] b,
    input     cin,
    output   cout,
    output [3:0] sum );
    
// Instantiate 100 copies of bcd_fadd to create a 100-digit BCD ripple-carry adder. 
//Your adder should add two 100-digit BCD numbers (packed into 400-bit vectors) 
//and a carry-in to produce a 100-digit sum and carry out.


// Hint: An instance array or generate statement would be useful here.

module top_module( 
    input [399:0] a, b,
    input cin,
    output cout,
    output [399:0] sum );
genvarii;
generatefor(ii=0;ii<100;ii=ii+1)
begin : bcd_fadd_gen
    wire [3:0] a_slice, b_slice, sum_slice;
    wire cout_slice;
    assign a_slice = a[ii*4+:4];
    assign b_slice = b[ii*4+:4];
    assign sum[ii*4+:4] = sum_slice;
    bcd_fadd u_bcd_fadd (
        .a(a_slice),
        .b(b_slice),
        .cin((ii == 0) ? cin : cout_slice),
        .cout((ii == 99) ? cout : cout_slice),
        .sum(sum_slice)
    );
end
endgenerate
endmodule