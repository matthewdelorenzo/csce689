    assign out = a & b;
endmodule
