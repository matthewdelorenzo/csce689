//Design a 16-bit adder.
//There are two 16 bit inputs (in1 and in2) and a single carry-in input bit, cin.
//The outputs are a 16 bit value, [15:0] sum, and a single carry-out output bit, cout.
//The module should utilize the inputs (in1 and in2) and the cin bit to obtain the output sum and cout values.
module top_module(output [15:0] sum,
                      output cout,
                      input [15:0] in1, in2,
                      input cin);
\n   assign sum = in1 + in2 + cin;\n  assign cout =(in1+in2 + cin) > 16'hFFFF;\nendmodule